-- Push Button Filter Module
-- This module implements debouncing filters for push button inputs
-- It uses a 4-bit shift register for each input to filter out noise and bounce
-------------------------------------------------------------------------------

-- Session 202, Team number 7, Bill Lu, Ailu Lin
library ieee;
use ieee.std_logic_1164.all;

entity PB_filters is port (
	-- Clock input for synchronization
	clkin				: in std_logic;
	-- Active-low reset input
	rst_n				: in std_logic;
	-- Filtered active-low reset output
	rst_n_filtered	: out std_logic;
	-- Active-low push button inputs
	pb_n				: in  std_logic_vector (3 downto 0);
	-- Filtered active-low push button outputs
	pb_n_filtered	: out	std_logic_vector(3 downto 0)							 
	); 
end PB_filters;

architecture ckt of PB_filters is

	-- Shift registers for debouncing each input
	-- sreg4: reset button
	-- sreg3-sreg0: push buttons 3-0
	Signal sreg0, sreg1, sreg2, sreg3, sreg4	: std_logic_vector(3 downto 0);

BEGIN

	-- Process to handle input filtering
	process (clkin) is

	begin
		if (rising_edge(clkin)) then
		
			-- Shift in new input values into shift registers
			-- Reset button shift register
			sreg4(3 downto 0) <= sreg4(2 downto 0) & rst_n;
				
			-- Push button shift registers
			sreg3(3 downto 0) <= sreg3(2 downto 0) & pb_n(3);
			sreg2(3 downto 0) <= sreg2(2 downto 0) & pb_n(2);
			sreg1(3 downto 0) <= sreg1(2 downto 0) & pb_n(1);
			sreg0(3 downto 0) <= sreg0(2 downto 0) & pb_n(0);
				
		end if;
		
		-- Generate filtered outputs using majority voting
		-- Output is 1 if at least 3 of the last 4 samples were 1
		rst_n_filtered   <= sreg4(3) OR sreg4(2) OR sreg4(1);
		
		pb_n_filtered(3) <= sreg3(3) OR sreg3(2) OR sreg3(1);
		pb_n_filtered(2) <= sreg2(3) OR sreg2(2) OR sreg2(1);
		pb_n_filtered(1) <= sreg1(3) OR sreg1(2) OR sreg1(1);
		pb_n_filtered(0) <= sreg0(3) OR sreg0(2) OR sreg0(1);
		
	end process;
end ckt;
